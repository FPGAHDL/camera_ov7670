module address_translator(h,v,address);

input [9:0] h;
input [9:0] v;
output [15:0] address;



endmodule
